/*
	Title: MIPS Single Cycle CPU Testbench
	Author: Selene (Computer System and Architecture Lab, ICE, CYCU) 
*/
module tb_SingleCycle ();
    reg clk, rst;

    // ���ͮɯߡA�g���G10ns
    initial begin
        clk = 1;
        forever #5 clk = ~clk;
    end

    initial begin
        $dumpfile("tb_SingleCycle.vcd");
        $dumpvars(3, CPU);
        #500;
        $finish;
        $stop();
    end


    initial begin
        rst = 1'b1;
        /*
			���O��ưO����A�ɦW"instr_mem.txt, data_mem.txt"�i�ۦ�ק�
			�C�@�欰1 Byte��ơA�H��Ӣ̤��i��Ʀr���
			�B��Little Endian�s�X
		*/
        $readmemh("instr_mem.txt", CPU.InstrMem.mem_array);
        $readmemh("data_mem.txt", CPU.DatMem.mem_array);
        // �]�w�Ȧs����l�ȡA�C�@�欰�@���Ȧs�����
        $readmemh("reg.txt", CPU.RegFile.file_array);
        #10;
        rst = 1'b0;
    end

    always @(posedge clk) begin
        $display("%d, PC:", $time / 10 - 1, CPU.pc);
        if (CPU.opcode == 6'd0) begin
            $display("%d, wd: %d", $time / 10 - 1, CPU.rfile_wd);
            if (CPU.funct == 6'd32) $display("%d, ADD\n", $time / 10 - 1);
            else if (CPU.funct == 6'd34) $display("%d, SUB\n", $time / 10 - 1);
            else if (CPU.funct == 6'd36) $display("%d, AND\n", $time / 10 - 1);
            else if (CPU.funct == 6'd37) $display("%d, OR\n", $time / 10 - 1);
        end else if (CPU.opcode == 6'd35) $display("%d, LW\n", $time / 10 - 1);
        else if (CPU.opcode == 6'd43) $display("%d, SW\n", $time / 10 - 1);
        else if (CPU.opcode == 6'd4) $display("%d, BEQ\n", $time / 10 - 1);
        else if (CPU.opcode == 6'd2) $display("%d, J\n", $time / 10 - 1);
    end

    mips_single CPU (
        clk,
        rst
    );

endmodule
